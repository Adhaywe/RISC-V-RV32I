//******************************************************************************************
// Design: mmu_wrapper.sv
// Author:
// Description: wrapper module that connects the mmu unit with the memory
// v 0.1
//******************************************************************************************
import types::*;

module mac_wrapper
(
    input  mac_op_t     mac_op,

    input  logic [31:0] mem_data1_i,    // matrix A elements from memory
    input  logic [31:0] mem_data2_i,
    input  logic [31:0] mem_data3_i,

    input  logic [31:0] mem_data4_i,    // matrix B elements from memory
    input  logic [31:0] mem_data5_i,
    input  logic [31:0] mem_data6_i,

    output logic [31:0] mem_data1_o,    // computed output to memory
    output logic [31:0] mem_data2_o,
    output logic [31:0] mem_data3_o
);

    logic [71:0] matA_i, matB_i;
    logic [71:0] res_o;


    assign matA_i = {mem_data1_i[7:0], mem_data1_i[15:8], mem_data1_i[23:16],
                     mem_data2_i[7:0], mem_data2_i[15:8], mem_data2_i[23:16],
                     mem_data3_i[7:0], mem_data3_i[15:8], mem_data3_i[23:16]};


    assign matB_i = {mem_data1_i[7:0], mem_data1_i[15:8], mem_data1_i[23:16],
                     mem_data2_i[7:0], mem_data2_i[15:8], mem_data2_i[23:16],
                     mem_data3_i[7:0], mem_data3_i[15:8], mem_data3_i[23:16]};


    mac mac_instance
    (
        .matrixA_i ( matA_i   ),
        .matrixB_i ( matB_i   ),
        .mac_op    ( mac_op   ),
        .result_o  ( res_o    )
    );

    assign mem_data1_o = {8'b0, res_o[71:64], res_o[63:56], res_o[55:48]};
    assign mem_data2_o = {8'b0, res_o[47:40], res_o[39:32], res_o[31:24]};
    assign mem_data3_o = {8'b0, res_o[23:16], res_o[15:8],  res_o[7:0]};

endmodule
