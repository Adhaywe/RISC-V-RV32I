//******************************************************************************************
// Design: adder.sv
// Author: Adam 
// Description: adder
// v 0.1
//******************************************************************************************


module adder (
	    input [31:0]  a, b,
		output [31:0] y
);

    assign y = a + b;

endmodule