package mac_pkg;

    localparam DATA_WIDTH = 72;
    localparam MAT_SIZE   = 3;
    localparam VAR_WIDTH  = 8;
    localparam MADD = 2'b00;
    localparam MSUB = 2'b01;
    localparam MMUL = 2'b10;

endpackage