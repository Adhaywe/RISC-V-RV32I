package mac_pkg;
    localparam DATA_WIDTH = 72;
    localparam MAT_SIZE   = 3;
    localparam VAR_WIDTH  = 8;

    localparam ADD = 2'b00;
    localparam SUB = 2'b01;
    localparam MUL = 2'b10;
    localparam MMUL = 2'b11;

endpackage